module Core(
    input clk,
    input reset
);

endmodule:Core