module Execute(
    //stage info
    id_stage.i id_info,
    ex_stage.o ex_info
);


endmodule