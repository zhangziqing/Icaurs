`define RESET_VECTOR 32'h01c000000