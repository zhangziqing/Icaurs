//basic width
`define DATA_WIDTH 32
`define ADDR_WIDTH 32
`define INST_WITDH 32
`define REG_WIDTH 5
`define REG_NUM 32

`define NUM_OF_BYTES 4


//implentation specific width

`define EXU_OP_WIDTH 6
`define EXU_OP_NUM 16


`define LSU_OP_WIDTH 4
`define LSU_OP_NUM 16