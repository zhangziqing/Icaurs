`define CSR_CRMD      14'h0
`define CSR_PRMD      14'h1
`define CSR_EUEN      14'h2
`define CSR_ECFG      14'h4
`define CSR_ESTAT     14'h5
`define CSR_ERA       14'h6
`define CSR_BADV      14'h7
`define CSR_EENTRY    14'hc
`define CSR_TLBIDX    14'h10
`define CSR_TLBEHI    14'h11
`define CSR_TLBELO0   14'h12
`define CSR_TLBELO1   14'h13
`define CSR_ASID      14'h18
`define CSR_PGDL      14'h19
`define CSR_PGDH      14'h1a
`define CSR_PGD       14'h1b
`define CSR_CPUID     14'h20
`define CSR_SAVE0     14'h30
`define CSR_SAVE1     14'h31
`define CSR_SAVE2     14'h32
`define CSR_SAVE3     14'h33
`define CSR_TID       14'h40
`define CSR_TCFG      14'h41
`define CSR_TVAL      14'h42
`define CSR_TICLR     14'h44
`define CSR_LLBCTL    14'h60
`define CSR_TLBRENTRY 14'h88
`define CSR_CTAG      14'h98
`define CSR_DMW0      14'h180
`define CSR_DMW1      14'h181
