module MemoryAccess(

);

endmodule:MemoryAccess