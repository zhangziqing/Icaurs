module BTB(
    
);


endmodule