module InstFecth(
    output  [`ADDR_WIDTH - 1 : 0 ]   pc,
    branch_info.i branch_info,
)

endmodule:InstFecth