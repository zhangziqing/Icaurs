`define ALU_OP_WIDTH 5
`define ALU_ADD 5'b00000
`define ALU_SUB 5'b00010
