module MemoryAccess(

);

endmodule:MemoryAccess