module InstCache(
    axi4_if.m axi4
);

endmodule