interface if_stage_if;



endinterface
