module Core(

);

endmodule:core