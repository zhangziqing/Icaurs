interface if_stage;



endinterface