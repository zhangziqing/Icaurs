`define CSR_CRMD      0x0
`define CSR_PRMD      0x1
`define CSR_EUEN      0x2
`define CSR_ECFG      0x4
`define CSR_ESTAT     0x5
`define CSR_ERA       0x6
`define CSR_BADV      0x7
`define CSR_EENTRY    0xc
`define CSR_TLBIDX    0x10
`define CSR_TLBEHI    0x11
`define CSR_TLBELO0   0x12
`define CSR_TLBELO1   0x13
`define CSR_ASID      0x18
`define CSR_PGDL      0x19
`define CSR_PGDH      0x1a
`define CSR_PGD       0x1b
`define CSR_CPUID     0x20
`define CSR_SAVE0     0x30
`define CSR_SAVE1     0x31
`define CSR_SAVE2     0x32
`define CSR_SAVE3     0x33
`define CSR_TID       0x40
`define CSR_TCFG      0x41
`define CSR_TVAL      0x42
`define CSR_TICLR     0x44
`define CSR_LLBCTL    0x60
`define CSR_TLBRENTRY 0x88
`define CSR_CTAG      0x98
`define CSR_DMW0      0x180
`define CSR_DMW1      0x181
